/media/emilio/Datos/Dropbox/Seven/IRIG-B/freq_div.vhd