LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY wb_irig_b IS
	GENERIC(
		FREQ_IN 		: IN		INTEGER:=62500000
	);
	PORT(    
		rst_n_i		: IN     STD_LOGIC;
		clk_sys_i	: IN     STD_LOGIC;
		wb_adr_i    : IN     STD_LOGIC_VECTOR(3 DOWNTO 0);
		wb_dat_i    : IN     STD_LOGIC_VECTOR(31 DOWNTO 0);
		wb_dat_o    : OUT    STD_LOGIC_VECTOR(31 DOWNTO 0);
		wb_cyc_i    : IN     STD_LOGIC;
		wb_sel_i    : IN     STD_LOGIC_VECTOR(3 DOWNTO 0);
		wb_stb_i    : IN     STD_LOGIC;
		wb_we_i     : IN     STD_LOGIC;
		wb_ack_o    : OUT    STD_LOGIC;
		wb_stall_o  : OUT    STD_LOGIC;
		wb_int_o    : OUT    STD_LOGIC;
		
		pps_in		: IN 		STD_LOGIC;
		output		: OUT 	STD_LOGIC
	);
END ENTITY wb_irig_b;


ARCHITECTURE funcional OF wb_irig_b IS
	COMPONENT irig_b
		GENERIC(
			FREQ_IN	:INTEGER := FREQ_IN
		);
	PORT(
		clk,reset,pps,enable,update	:IN STD_LOGIC;
		output			:OUT STD_LOGIC;
		irq_ou			:OUT STD_LOGIC;
		year				:IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		day				:IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		hour				:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		min				:IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		sec				:IN STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
	END COMPONENT;
	COMPONENT wb_irigb
	PORT(
		rst_n_i                                  : IN     STD_LOGIC;
		clk_sys_i                                : IN     STD_LOGIC;
		wb_adr_i                                 : IN     STD_LOGIC_vector(3 downto 0);
		wb_dat_i                                 : IN     STD_LOGIC_vector(31 downto 0);
		wb_dat_o                                 : OUT    STD_LOGIC_vector(31 downto 0);
		wb_cyc_i                                 : IN     STD_LOGIC;
		wb_sel_i                                 : IN     STD_LOGIC_vector(3 downto 0);
		wb_stb_i                                 : IN     STD_LOGIC;
		wb_we_i                                  : IN     STD_LOGIC;
		wb_ack_o                                 : OUT    STD_LOGIC;
		wb_stall_o                               : OUT    STD_LOGIC;
		wb_int_o                                 : OUT    STD_LOGIC;
	
		irigb_stat_res_o                         : OUT    STD_LOGIC;
		irigb_stat_ena_o                         : OUT    STD_LOGIC;
		irigb_yea_year_o                         : OUT    STD_LOGIC_VECTOR(31 downto 0);
		irigb_day_day_o                          : OUT    STD_LOGIC_VECTOR(31 downto 0);
		irigb_hou_hou_o                          : OUT    STD_LOGIC_VECTOR(31 downto 0);
		irigb_min_min_o                          : OUT    STD_LOGIC_VECTOR(31 downto 0);
		irigb_sec_sec_o                          : OUT    STD_LOGIC_VECTOR(31 downto 0);
		irq_hur_i                                : IN     STD_LOGIC
	);
	END COMPONENT;
	SIGNAL rst_prev,up,rs				: STD_LOGIC:='0';
	
	SIGNAL year,day,hour,min,sec		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL irq,res,en						: STD_LOGIC;
BEGIN
	irig: irig_b
		GENERIC MAP(
			FREQ_IN
		)
		PORT MAP(
			clk_sys_i,
			res,
			pps_in,
			en,
			up,
			output,
			irq,
			year(11 DOWNTO 0),
			day(8 DOWNTO 0),
			hour(4 DOWNTO 0),
			min(5 DOWNTO 0),
			sec(5 DOWNTO 0)
		);
	wb_if: wb_irigb
		PORT MAP(
			rst_n_i,
			clk_sys_i,
			wb_adr_i,
			wb_dat_i,
			wb_dat_o,
			wb_cyc_i,
			wb_sel_i,
			wb_stb_i,
			wb_we_i,
			wb_ack_o,
			wb_stall_o,
			wb_int_o,
			rs,
			en,
			year,
			day,
			hour,
			min,
			sec,
			irq
		);
	
	PROCESS(clk_sys_i)
	BEGIN
		IF rising_edge(clk_sys_i) THEN
			IF(wb_we_i='1') and (wb_adr_i/="0000")THEN
				up<='1';
			ELSE
				up<='0';
			END IF;
		END IF;
	END PROCESS;
	
	
	ctrlrst: PROCESS(clk_sys_i)
	BEGIN
		IF rising_edge(clk_sys_i) THEN
			rst_prev<=rs;
		END IF;
	END PROCESS ctrlrst;
	
	res<='1' WHEN (rst_n_i='0') or (rst_prev='0' and res='1') ELSE '0';
END ARCHITECTURE funcional;

















