/media/emilio/Datos/Dropbox/Seven/IRIG-B/irigb_mod.vhd