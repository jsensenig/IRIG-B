/media/emilio/Datos/Dropbox/Seven/IRIG-B/irig_b.vhd